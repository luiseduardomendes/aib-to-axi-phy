// ============================================================================
// Description: Top-Level Wrapper for the AIB to AXI Integrated System
//
// Purpose:
// This module wraps the entire 'aib_axi_top' system. It provides a clean
// instantiation point for integrating the complete leader/follower bridge
// system into a larger design, such as a full SoC or testbench.
//
// Instantiates:
// 1. aib_axi_m2s2_top (Corrected name from comments)
// ============================================================================

module aib_axi_top_wrapper #(
    // --- Parameters are passed directly to the core aib_axi_top module ---
    parameter ACTIVE_CHNLS      = 1,
    parameter NBR_CHNLS         = 24,
    parameter LEADER_NBR_BUMPS  = 102,
    parameter FOLLOWER_NBR_BUMPS= 102,
    parameter NBR_PHASES        = 4,
    parameter NBR_LANES         = 40,
    parameter MS_SSR_LEN        = 81,
    parameter SL_SSR_LEN        = 73,
    parameter DWIDTH            = 40,
    parameter AXI_CHNL_NUM      = 1,
    parameter ADDRWIDTH         = 32,
    parameter IDWIDTH           = 4,
    parameter GEN2_MODE         = 1'b1
) (
    // ========================================================================
    // Leader (Master Bridge) Interface
    // ========================================================================
    inout leader_vddc1,
    inout leader_vddc2,
    inout leader_vddtx,
    inout leader_vss,
    input   leader_m_wr_clk,
    input   leader_m_rd_clk,
    input   leader_m_fwd_clk,
    input leader_i_osc_clk,
    input  [NBR_CHNLS-1: 0] leader_ns_adapter_rstn,
    input  [NBR_CHNLS-1: 0] leader_ns_mac_rdy,
    output [NBR_CHNLS-1: 0] leader_fs_mac_rdy,
    output [NBR_CHNLS-1: 0] leader_m_rx_align_done,
    input leader_avmm_clk,
    input leader_avmm_rst_n,
    input leader_i_cfg_avmm_clk,
    input leader_i_cfg_avmm_rst_n,
    input [16:0] leader_i_cfg_avmm_addr,
    input [3:0] leader_i_cfg_avmm_byte_en,
    input leader_i_cfg_avmm_read,
    input leader_i_cfg_avmm_write,
    input [31:0] leader_i_cfg_avmm_wdata,
    output leader_o_cfg_avmm_rdatavld,
    output [31:0] leader_o_cfg_avmm_rdata,
    output leader_o_cfg_avmm_waitreq,
    input leader_clk_wr,
    input leader_rst_wr_n,
    // CORRECTED CREDITS: Leader (AXI Slave) needs R and B credits
    input [7:0] follower_init_r_credit,
    input [7:0] follower_init_b_credit,
    input [15:0] leader_delay_x_value,
    input [15:0] leader_delay_y_value,
    input [15:0] leader_delay_z_value,
    input  [IDWIDTH-1:0]     s_axi_awid,
    input  [ADDRWIDTH-1:0]   s_axi_awaddr,
    input  [7:0]             s_axi_awlen,
    input  [2:0]             s_axi_awsize,
    input  [1:0]             s_axi_awburst,
    input                    s_axi_awvalid,
    output                   s_axi_awready,
    input  [IDWIDTH-1:0]     s_axi_wid,
    input  [127:0]           s_axi_wdata,
    input  [15:0]            s_axi_wstrb,
    input                    s_axi_wlast,
    input                    s_axi_wvalid,
    output                   s_axi_wready,
    output [IDWIDTH-1:0]     s_axi_bid,
    output [1:0]             s_axi_bresp,
    output                   s_axi_bvalid,
    input                    s_axi_bready,
    input  [IDWIDTH-1:0]     s_axi_arid,
    input  [ADDRWIDTH-1:0]   s_axi_araddr,
    input  [7:0]             s_axi_arlen,
    input  [2:0]             s_axi_arsize,
    input  [1:0]             s_axi_arburst,
    input                    s_axi_arvalid,
    output                   s_axi_arready,
    output [IDWIDTH-1:0]     s_axi_rid,
    output [127:0]           s_axi_rdata,
    output [1:0]             s_axi_rresp,
    output                   s_axi_rlast,
    output                   s_axi_rvalid,
    input                    s_axi_rready,

    // ========================================================================
    // Follower (Slave Bridge) Interface
    // ========================================================================
    inout follower_vddc1,
    inout follower_vddc2,
    inout follower_vddtx,
    inout follower_vss,
    input   follower_m_wr_clk,
    input   follower_m_rd_clk,
    input   follower_m_fwd_clk,
    input  [NBR_CHNLS-1: 0] follower_ns_adapter_rstn,
    input  [NBR_CHNLS-1: 0] follower_ns_mac_rdy,
    output [NBR_CHNLS-1: 0] follower_fs_mac_rdy,
    output [NBR_CHNLS-1: 0] follower_m_rx_align_done,
    output [NBR_CHNLS-1: 0] follower_ms_tx_transfer_en,
    output [NBR_CHNLS-1: 0] follower_sl_tx_transfer_en,
    input  follower_clk_wr,
    input  follower_rst_wr_n,
    // CORRECTED CREDITS: Follower (AXI Master) needs AR, AW, and W credits
    input [7:0] leader_init_ar_credit,
    input [7:0] leader_init_aw_credit,
    input [7:0] leader_init_w_credit,
    input [15:0] follower_delay_x_value,
    input [15:0] follower_delay_y_value,
    input [15:0] follower_delay_z_value,
    // --- Follower Avalon MM Interface ---
    input  follower_avmm_clk,
    input  follower_avmm_rst_n,
    input  follower_i_cfg_avmm_clk,
    input  follower_i_cfg_avmm_rst_n,
    input  [16:0] follower_i_cfg_avmm_addr,
    input  [3:0]  follower_i_cfg_avmm_byte_en,
    input         follower_i_cfg_avmm_read,
    input         follower_i_cfg_avmm_write,
    input  [31:0] follower_i_cfg_avmm_wdata,
    output        follower_o_cfg_avmm_rdatavld,
    output [31:0] follower_o_cfg_avmm_rdata,
    output        follower_o_cfg_avmm_waitreq,
    output [IDWIDTH-1:0]     m_axi_awid,
    output [ADDRWIDTH-1:0]   m_axi_awaddr,
    output [7:0]             m_axi_awlen,
    output [2:0]             m_axi_awsize,
    output [1:0]             m_axi_awburst,
    output                   m_axi_awvalid,
    input                    m_axi_awready,
    output [IDWIDTH-1:0]     m_axi_wid,
    output [127:0]           m_axi_wdata,
    output [15:0]            m_axi_wstrb,
    output                   m_axi_wlast,
    output                   m_axi_wvalid,
    input                    m_axi_wready,
    input  [IDWIDTH-1:0]     m_axi_bid,
    input  [1:0]             m_axi_bresp,
    input                    m_axi_bvalid,
    output                   m_axi_bready,
    output [IDWIDTH-1:0]     m_axi_arid,
    output [ADDRWIDTH-1:0]   m_axi_araddr,
    output [7:0]             m_axi_arlen,
    output [2:0]             m_axi_arsize,
    output [1:0]             m_axi_arburst,
    output                   m_axi_arvalid,
    input                    m_axi_arready,
    input  [IDWIDTH-1:0]     m_axi_rid,
    input  [127:0]           m_axi_rdata,
    input  [1:0]             m_axi_rresp,
    input                    m_axi_rlast,
    input                    m_axi_rvalid,
    output                   m_axi_rready
);

    // ============================================================================
    // Core AIB AXI System Instantiation
    // ============================================================================
    aib_axi_m2s2_top #(
        .ACTIVE_CHNLS    (ACTIVE_CHNLS),
        .NBR_CHNLS       (NBR_CHNLS),
        .LEADER_NBR_BUMPS  (LEADER_NBR_BUMPS),
        .FOLLOWER_NBR_BUMPS(FOLLOWER_NBR_BUMPS),
        .NBR_PHASES      (NBR_PHASES),
        .NBR_LANES       (NBR_LANES),
        .MS_SSR_LEN      (MS_SSR_LEN),
        .SL_SSR_LEN      (SL_SSR_LEN),
        .DWIDTH          (DWIDTH),
        .AXI_CHNL_NUM    (AXI_CHNL_NUM),
        .ADDRWIDTH       (ADDRWIDTH),
        .IDWIDTH         (IDWIDTH),
        .GEN2_MODE       (GEN2_MODE)
    )
    u_aib_axi_top (
        // --- Leader Interface Connections ---
        .leader_vddc1(leader_vddc1),
        .leader_vddc2(leader_vddc2),
        .leader_vddtx(leader_vddtx),
        .leader_vss(leader_vss),
        .leader_m_wr_clk(leader_m_wr_clk),
        .leader_m_rd_clk(leader_m_rd_clk),
        .leader_m_fwd_clk(leader_m_fwd_clk),
        .leader_i_osc_clk(leader_i_osc_clk),
        .leader_ns_adapter_rstn(leader_ns_adapter_rstn),
        .leader_ns_mac_rdy(leader_ns_mac_rdy),
        .leader_fs_mac_rdy(leader_fs_mac_rdy),
        .leader_m_rx_align_done(leader_m_rx_align_done),
        .leader_avmm_clk(leader_avmm_clk),
        .leader_avmm_rst_n(leader_avmm_rst_n),
        .leader_i_cfg_avmm_clk(leader_i_cfg_avmm_clk),
        .leader_i_cfg_avmm_rst_n(leader_i_cfg_avmm_rst_n),
        .leader_i_cfg_avmm_addr(leader_i_cfg_avmm_addr),
        .leader_i_cfg_avmm_byte_en(leader_i_cfg_avmm_byte_en),
        .leader_i_cfg_avmm_read(leader_i_cfg_avmm_read),
        .leader_i_cfg_avmm_write(leader_i_cfg_avmm_write),
        .leader_i_cfg_avmm_wdata(leader_i_cfg_avmm_wdata),
        .leader_o_cfg_avmm_rdatavld(leader_o_cfg_avmm_rdatavld),
        .leader_o_cfg_avmm_rdata(leader_o_cfg_avmm_rdata),
        .leader_o_cfg_avmm_waitreq(leader_o_cfg_avmm_waitreq),
        .leader_clk_wr(leader_clk_wr),
        .leader_rst_wr_n(leader_rst_wr_n),
        .leader_init_ar_credit(leader_init_ar_credit),
        .leader_init_aw_credit(leader_init_aw_credit),
        .leader_init_w_credit(leader_init_w_credit),
        .leader_delay_x_value(leader_delay_x_value),
        .leader_delay_y_value(leader_delay_y_value),
        .leader_delay_z_value(leader_delay_z_value),
        .s_axi_awid(s_axi_awid),
        .s_axi_awaddr(s_axi_awaddr),
        .s_axi_awlen(s_axi_awlen),
        .s_axi_awsize(s_axi_awsize),
        .s_axi_awburst(s_axi_awburst),
        .s_axi_awvalid(s_axi_awvalid),
        .s_axi_awready(s_axi_awready),
        .s_axi_wid(s_axi_wid),
        .s_axi_wdata(s_axi_wdata),
        .s_axi_wstrb(s_axi_wstrb),
        .s_axi_wlast(s_axi_wlast),
        .s_axi_wvalid(s_axi_wvalid),
        .s_axi_wready(s_axi_wready),
        .s_axi_bid(s_axi_bid),
        .s_axi_bresp(s_axi_bresp),
        .s_axi_bvalid(s_axi_bvalid),
        .s_axi_bready(s_axi_bready),
        .s_axi_arid(s_axi_arid),
        .s_axi_araddr(s_axi_araddr),
        .s_axi_arlen(s_axi_arlen),
        .s_axi_arsize(s_axi_arsize),
        .s_axi_arburst(s_axi_arburst),
        .s_axi_arvalid(s_axi_arvalid),
        .s_axi_arready(s_axi_arready),
        .s_axi_rid(s_axi_rid),
        .s_axi_rdata(s_axi_rdata),
        .s_axi_rresp(s_axi_rresp),
        .s_axi_rlast(s_axi_rlast),
        .s_axi_rvalid(s_axi_rvalid),
        .s_axi_rready(s_axi_rready),

        // --- Follower Interface Connections ---
        .follower_vddc1(follower_vddc1),
        .follower_vddc2(follower_vddc2),
        .follower_vddtx(follower_vddtx),
        .follower_vss(follower_vss),
        .follower_m_wr_clk(follower_m_wr_clk),
        .follower_m_rd_clk(follower_m_rd_clk),
        .follower_m_fwd_clk(follower_m_fwd_clk),
        .follower_ns_adapter_rstn(follower_ns_adapter_rstn),
        .follower_ns_mac_rdy(follower_ns_mac_rdy),
        .follower_fs_mac_rdy(follower_fs_mac_rdy),
        .follower_m_rx_align_done(follower_m_rx_align_done),
        .follower_ms_tx_transfer_en(follower_ms_tx_transfer_en),
        .follower_sl_tx_transfer_en(follower_sl_tx_transfer_en),
        .follower_clk_wr(follower_clk_wr),
        .follower_rst_wr_n(follower_rst_wr_n),
        // CORRECTED CREDIT CONNECTIONS
        .follower_init_r_credit(follower_init_r_credit),
        .follower_init_b_credit(follower_init_b_credit),
        .follower_delay_x_value(follower_delay_x_value),
        .follower_delay_y_value(follower_delay_y_value),
        .follower_delay_z_value(follower_delay_z_value),
        // Avalon MM Interface
        .follower_avmm_clk(follower_avmm_clk),
        .follower_avmm_rst_n(follower_avmm_rst_n),
        .follower_i_cfg_avmm_clk(follower_i_cfg_avmm_clk),
        .follower_i_cfg_avmm_rst_n(follower_i_cfg_avmm_rst_n),
        .follower_i_cfg_avmm_addr(follower_i_cfg_avmm_addr),
        .follower_i_cfg_avmm_byte_en(follower_i_cfg_avmm_byte_en),
        .follower_i_cfg_avmm_read(follower_i_cfg_avmm_read),
        .follower_i_cfg_avmm_write(follower_i_cfg_avmm_write),
        .follower_i_cfg_avmm_wdata(follower_i_cfg_avmm_wdata),
        .follower_o_cfg_avmm_rdatavld(follower_o_cfg_avmm_rdatavld),
        .follower_o_cfg_avmm_rdata(follower_o_cfg_avmm_rdata),
        .follower_o_cfg_avmm_waitreq(follower_o_cfg_avmm_waitreq),
        .m_axi_awid(m_axi_awid),
        .m_axi_awaddr(m_axi_awaddr),
        .m_axi_awlen(m_axi_awlen),
        .m_axi_awsize(m_axi_awsize),
        .m_axi_awburst(m_axi_awburst),
        .m_axi_awvalid(m_axi_awvalid),
        .m_axi_awready(m_axi_awready),
        .m_axi_wid(m_axi_wid),
        .m_axi_wdata(m_axi_wdata),
        .m_axi_wstrb(m_axi_wstrb),
        .m_axi_wlast(m_axi_wlast),
        .m_axi_wvalid(m_axi_wvalid),
        .m_axi_wready(m_axi_wready),
        .m_axi_bid(m_axi_bid),
        .m_axi_bresp(m_axi_bresp),
        .m_axi_bvalid(m_axi_bvalid),
        .m_axi_bready(m_axi_bready),
        .m_axi_arid(m_axi_arid),
        .m_axi_araddr(m_axi_araddr),
        .m_axi_arlen(m_axi_arlen),
        .m_axi_arsize(m_axi_arsize),
        .m_axi_arburst(m_axi_arburst),
        .m_axi_arvalid(m_axi_arvalid),
        .m_axi_arready(m_axi_arready),
        .m_axi_rid(m_axi_rid),
        .m_axi_rdata(m_axi_rdata),
        .m_axi_rresp(m_axi_rresp),
        .m_axi_rlast(m_axi_rlast),
        .m_axi_rvalid(m_axi_rvalid),
        .m_axi_rready(m_axi_rready)
    );

endmodule